module routes

pub struct Router {
pub:
	route_name string
}
