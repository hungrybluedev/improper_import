module main

import app

fn main() {
	mut app := app.new_app()!
	app.run()
}
